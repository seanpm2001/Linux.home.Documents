-- Start of script
-- I have chosen VHDL as the 5th project language file for this project (WacOS) as along with Assembly, it is needed for hardware virtualization.
-- File version: 1 (Tuesday, April 27th 2021 at 8:00 pm)
-- File type: Virtual Hard Disk Language (VHDL) Source file (*.vhdl, *.vhd, *.vdi)
-- Line count (including blank lines and compiler line): 7
-- End of script

